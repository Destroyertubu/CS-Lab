`timescale 1ns/1ps

module AND(input A, input B, output out);

    assign out = A & B;
    
endmodule